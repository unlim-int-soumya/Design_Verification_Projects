import uvm_pkg::*;
`include "uvm_macros.svh"


`include "transaction.sv"
`include "generator.sv"
`include "driver.sv"
`include "monitor.sv"

`include "ref_model.sv"
`include "scoreboard.sv"
`include "agent.sv"
`include "env.sv"
`include "test.sv"