//package apb_pkg;
`include "apb_common.sv"
`include "apb_txn.sv"
`include "apb_gen.sv"
`include "apb_bfm.sv"
`include "apb_mon.sv"
`include "apb_agent.sv"
`include "apb_scb.sv"
`include "apb_cov_collecter.sv"
`include "apb_env.sv"
//endpackage
