program apb_base_test();
  apb_env env;
  
  initial begin
    env = new();
    env.run();
  end
  
endprogram
