
`ifndef IN_LENGTH
`define IN_LENGTH 16
`endif

`ifndef SEL_LENGTH
`define SEL_LENGTH 4
`endif

module mux_16x1(
  input [`SEL_LENGTH-1:0] sel, 
  input [`IN_LENGTH-1:0]in,
  input rstn,
  output reg out
);
  
  always @ (*) begin
    if(!rstn) begin
      out = 0;
    end else begin
      case(sel)
       	4'b0000: out = in[0];
        4'b0001: out = in[1];
        4'b0010: out = in[2];
        4'b0011: out = in[3];
        4'b0100: out = in[4];
        4'b0101: out = in[5];
        4'b0110: out = in[6];
        4'b0111: out = in[7];
        4'b1000: out = in[8];
        4'b1001: out = in[9];
        4'b1010: out = in[10];
        4'b1011: out = in[11];
        4'b1100: out = in[12];
        4'b1101: out = in[13];
        4'b1110: out = in[14];
        4'b1111: out = in[15]; 
        default: out = 0; 
      endcase
 	 end
  end

endmodule
